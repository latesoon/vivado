`timescale 1ns / 1ps
module multiply(              // �˷���
    input         clk,        // ʱ��
    input         mult_begin, // �˷���ʼ�ź�
    input  [31:0] mult_op1,   // �˷�Դ������1
    input  [31:0] mult_op2,   // �˷�Դ������2
    output [63:0] product,    // �˻�
    output        mult_end    // �˷������ź�
);

    //�˷����������źźͽ����ź�
    reg mult_valid;
    assign mult_end = mult_valid & ~(|multiplier) & (op2_sign | ~(xmultiplier)) ; //�˷������źţ�����ȫ0
    always @(posedge clk)
    begin
        if (!mult_begin || mult_end)
        begin
            mult_valid <= 1'b0;
        end
        else
        begin
            mult_valid <= 1'b1;
        end
    end

    //����Դ����ȡ����ֵ�������ľ���ֵΪ�䱾�������ľ���ֵΪȡ����1
    wire        op1_sign;      //������1�ķ���λ
    wire        op2_sign;      //������2�ķ���λ
    wire [31:0] op1;  //������1�ľ���ֵ
    wire [31:0] op2;  //������2�ľ���ֵ
    assign op1_sign = mult_op1[31];
    assign op2_sign = mult_op2[31];
    assign op1=mult_op1;
    assign op2=mult_op2;

    //���ر�����������ʱÿ������һλ
    reg  [63:0] multiplicand;
    reg  [63:0] m_multiplicand;
    always @ (posedge clk)
    begin
        if (mult_valid)
        begin    // ������ڽ��г˷����򱻳���ÿʱ������һλ
            multiplicand <= {multiplicand[61:0],2'b0};
            m_multiplicand <= {m_multiplicand[61:0],2'b0};
        end
        else if (mult_begin) 
        begin   // �˷���ʼ�����ر�������Ϊ����1�ľ���ֵ
            if(op1_sign)
            begin
                multiplicand <= {32'hFFFF_FFFF,op1};
                m_multiplicand <={31'b0,(~op1+1),1'b0};
            end
            else
            begin
                multiplicand <= {32'b0,op1};
                m_multiplicand<= {31'h7FFF_FFFF,(~op1+1),1'b0};
            end
        end
    end

    //���س���������ʱÿ������һλ
    reg  [31:0] multiplier;
    reg  xmultiplier;
    always @ (posedge clk)
    begin
        if (mult_valid)
        begin   // ������ڽ��г˷��������ÿʱ������һλ
            xmultiplier <= multiplier[1];
            multiplier <= {2'b0,multiplier[31:2]}; 
        end
        else if (mult_begin)
        begin   // �˷���ʼ�����س�����Ϊ����2�ľ���ֵ
            multiplier <= op2;
            xmultiplier<= 1'b0;
        end
    end
    
    // ���ֻ�������ĩλΪ1���ɱ��������Ƶõ�������ĩλΪ0�����ֻ�Ϊ0
    wire [63:0] partial_product;
    assign partial_product = mult_end?64'b0:((xmultiplier ? multiplicand : 64'b0)+(multiplier[0] ? multiplicand: 64'b0)+(multiplier[1]?m_multiplicand:64'b0));
    
    //�ۼ���
    reg [63:0] product_temp;
    always @ (posedge clk)
    begin
        if (mult_valid)
        begin
            product_temp <= product_temp + partial_product;
        end
        else if (mult_begin) 
        begin
            product_temp <= 64'd0;  // �˷���ʼ���˻����� 
        end
    end 
    //���˷����Ϊ����������Ҫ�Խ��ȡ��+1
    assign product = product_temp;
endmodule
